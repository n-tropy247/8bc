* SN74LS04 Hex Inverter Simulation

* Define the power supply
VCC 14 0 DC 5V

* Define the ground
VSS 7 0 0V

* Define input signals for all inverters
V1 1 0 PULSE(0 5 0 10n 10n 20n 40n)  * Pulse signal for input 1A
V2 3 0 PULSE(0 5 10n 10n 10n 20n 40n) * Pulse signal for input 2A
V3 5 0 PULSE(0 5 20n 10n 10n 20n 40n) * Pulse signal for input 3A
V4 9 0 PULSE(0 5 30n 10n 10n 20n 40n) * Pulse signal for input 4A
V5 11 0 PULSE(0 5 40n 10n 10n 20n 40n) * Pulse signal for input 5A
V6 13 0 PULSE(0 5 50n 10n 10n 20n 40n) * Pulse signal for input 6A

* Inverter connections
X1 1 2 3 4 5 6 7 8 9 10 11 12 13 14 SN74LS04

* Subcircuit definition for SN74LS04 with all 14 pins
.subckt SN74LS04 1A 1Y 2A 2Y 3A 3Y GND 4Y 4A 5Y 5A 6Y 6A VCC
* Inverter 1
M1 1Y 1A VCC VCC PMOS L=1u W=1u
M2 1Y 1A GND GND NMOS L=1u W=1u
R1 1Y VCC 10k
* Inverter 2
M3 2Y 2A VCC VCC PMOS L=1u W=1u
M4 2Y 2A GND GND NMOS L=1u W=1u
R2 2Y VCC 10k
* Inverter 3
M5 3Y 3A VCC VCC PMOS L=1u W=1u
M6 3Y 3A GND GND NMOS L=1u W=1u
R3 3Y VCC 10k
* Inverter 4
M7 4Y 4A VCC VCC PMOS L=1u W=1u
M8 4Y 4A GND GND NMOS L=1u W=1u
R4 4Y VCC 10k
* Inverter 5
M9 5Y 5A VCC VCC PMOS L=1u W=1u
M10 5Y 5A GND GND NMOS L=1u W=1u
R5 5Y VCC 10k
* Inverter 6
M11 6Y 6A VCC VCC PMOS L=1u W=1u
M12 6Y 6A GND GND NMOS L=1u W=1u
R6 6Y VCC 10k
.ends SN74LS04

* Simulation control
.tran 0.1n 100n

* Outputs
.print tran V(2) V(4) V(6) V(8) V(10) V(12)

.end
